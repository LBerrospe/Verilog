`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Universidad de Gualadajara
// Engineer: Hector Eduardo Berrospe Barajas
// 
// Create Date: 13.05.2016 18:03:32
// Design Name: Decode
// Module Name: Decode
// Project Name: Processor
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Decoder(
        input [4:0] w_addr,
        input en_addr,
        output reg [31:0] out
    );
    
    always@*
    begin
        case(en_addr)
            1'b0: out = 32'b00000000000000000000000000000000;
            1'b1:
            begin
                case(w_addr)
                    5'b 00000: out = 32'b00000000000000000000000000000001;
                    5'b 00001: out = 32'b00000000000000000000000000000010;
                    5'b 00010: out = 32'b00000000000000000000000000000100;
                    5'b 00011: out = 32'b00000000000000000000000000001000;
                    5'b 00100: out = 32'b00000000000000000000000000010000;
                    5'b 00101: out = 32'b00000000000000000000000000100000;
                    5'b 00110: out = 32'b00000000000000000000000001000000;
                    5'b 00111: out = 32'b00000000000000000000000010000000;
                    5'b 01000: out = 32'b00000000000000000000000100000000;
                    5'b 01001: out = 32'b00000000000000000000001000000000;
                    5'b 01010: out = 32'b00000000000000000000010000000000;
                    5'b 01011: out = 32'b00000000000000000000100000000000;
                    5'b 01100: out = 32'b00000000000000000001000000000000;
                    5'b 01101: out = 32'b00000000000000000010000000000000;
                    5'b 01110: out = 32'b00000000000000000100000000000000;
                    5'b 01111: out = 32'b00000000000000001000000000000000;
                    5'b 10000: out = 32'b00000000000000010000000000000000;
                    5'b 10001: out = 32'b00000000000000100000000000000000;
                    5'b 10010: out = 32'b00000000000001000000000000000000;
                    5'b 10011: out = 32'b00000000000010000000000000000000;
                    5'b 10100: out = 32'b00000000000100000000000000000000;
                    5'b 10101: out = 32'b00000000001000000000000000000000;
                    5'b 10110: out = 32'b00000000010000000000000000000000;
                    5'b 10111: out = 32'b00000000100000000000000000000000;
                    5'b 11000: out = 32'b00000001000000000000000000000000;
                    5'b 11001: out = 32'b00000010000000000000000000000000;
                    5'b 11010: out = 32'b00000100000000000000000000000000;
                    5'b 11011: out = 32'b00001000000000000000000000000000;
                    5'b 11100: out = 32'b00010000000000000000000000000000;
                    5'b 11101: out = 32'b00100000000000000000000000000000;
                    5'b 11110: out = 32'b01000000000000000000000000000000;
                    5'b 11111: out = 32'b10000000000000000000000000000000;
                    
                    default: out = 32'b00000000000000000000000000000000;
                endcase
            end
            default: out = 32'b00000000000000000000000000000000;
        endcase
    end
endmodule
