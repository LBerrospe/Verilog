`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Universidad de Gualadajara
// Engineer: Hector Eduardo Berrospe Barajas
// 
// Create Date: 30.04.2016 21:24:48
// Design Name: ROM_I
// Module Name: ROM_I
// Project Name: Processor
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module ROM_I(
    input [3:0] addr_ROM,
    output reg [31:0] d
    );
    
    always@*
    begin
			case(addr_ROM)
				4'b0000 : d <=  32'b00000000010000010000000000000010;
				4'b0001 : d <=  32'b00000000001000100000000000000110; 
				4'b0010 : d <=  32'b00001000001000100000000000000010; 
				4'b0011 : d <=  32'b00000000000000000000000000000101;
				4'b0100 : d <=  32'b00000000000000000000000000000110;
				4'b0101 : d <=  32'b00000000000000000000000000000110; 
				4'b0110 : d <=  32'b00000000000000000000000000000111; 
				4'b0111 : d <=  32'b00000000000000000000000000001000; 
				4'b1000 : d <=  32'b00000000000000000000000000001001; 
				4'b1001 : d <=  32'b00000000000000000000000000001010; 
				4'b1010 : d <=  32'b00000000000000000000000000001011;
				4'b1011 : d <=  32'b00000000000000000000000000001100;
				4'b1100 : d <=  32'b00000000000000000000000000001101;
				4'b1101 : d <=  32'b00000000000000000000000000001110;
				4'b1110 : d <=  32'b00000000000000000000000000000000; 
                4'b1111 : d <=  32'b00000000000000000000000000000001; 

				default : d <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;	

		endcase//FIN case en          
    end
endmodule
