`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.04.2016 21:24:48
// Design Name: 
// Module Name: ROM_I
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module ROM_I(
    input [3:0] addr_ROM,
    output reg [31:0] d
    );
    
    always@*
    begin
			case(addr_ROM)
				4'b0000 : d <=  32'b00000000000000000000000000000100;
				4'b0001 : d <=  32'b00000000000000000000000000000100; 
				4'b0010 : d <=  32'b00000000000000000000000000000101;
				4'b0011 : d <=  32'b00000000000000000000000000000101;
				4'b0100 : d <=  32'b00000000000000000000000000000110;
				4'b0101 : d <=  32'b00000000000000000000000000000110; 
				4'b0110 : d <=  32'b00000000000000000000000000000111; 
				4'b0111 : d <=  32'b00000000000000000000000000001000; 
				4'b1000 : d <=  32'b00000000000000000000000000001001; 
				4'b1001 : d <=  32'b00000000000000000000000000001010; 
				4'b1010 : d <=  32'b00000000000000000000000000001011;
				4'b1011 : d <=  32'b00000000000000000000000000001100;
				4'b1100 : d <=  32'b00000000000000000000000000001101;
				4'b1101 : d <=  32'b00000000000000000000000000001110;
				4'b1110 : d <=  32'b00000000000000000000000000000000; //Lee arit
                4'b1111 : d <=  32'b00000000000000000000000000000001; //Lee Log  


				default : d <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;	

		endcase//FIN case en          
    end
endmodule
