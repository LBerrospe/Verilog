`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.04.2016 21:25:42
// Design Name: 
// Module Name: ROM_OP2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module ROM_OP2(
    input en_ROM,
    input [3:0] addr_ROM,
    output reg [31:0] d
    );
    
    always@*
    begin
		case(en_ROM)
		1'b1:
			case(addr_ROM)
                4'b0000 : d <=  32'b00000000000000000000000000000101; 
                4'b0001 : d <=  32'b00000000000000000000000000000111;
                4'b0010 : d <=  32'b00000000000000000000000000001110; 
                4'b0011 : d <=  32'b00000000000000000000000000001111; 
                4'b0100 : d <=  32'b00000000000000000000000000011111; 
                4'b0101 : d <=  32'b00000000000000000000000000110111; 
                4'b0110 : d <=  32'b00000000000000000000000001010111; 
                4'b0111 : d <=  32'b00000000000000000000000000111111;
                4'b1000 : d <=  32'b00000000000000000000000000110000;
                4'b1001 : d <=  32'b00000000000000000000000000110010;
                4'b1010 : d <=  32'b00000000000000000000000000110001;
                4'b1011 : d <=  32'b00000000000000000000000000110110;
                4'b1100 : d <=  32'b00000000000000000000000000101111;
                4'b1101 : d <=  32'b00000000000000000000000010010000;
                4'b1110 : d <=  32'b00000000000000000000000001101000;    
                4'b1111 : d <=  32'b00000000000000000000000001101001;    

				default : d <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;	
			endcase//FIN case addr
			
			default : d <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
		endcase//FIN case en          
    end
endmodule