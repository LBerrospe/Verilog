`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.04.2016 21:25:17
// Design Name: 
// Module Name: ROM_OP1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module ROM_OP1(
    input en_ROM,
    input [3:0] addr_ROM,
    output reg [31:0] d
    );
    
    always@*
    begin
		case(en_ROM)
		1'b1:
			case(addr_ROM)
				4'b0000 : d <=  32'b00000000000000000000000000000100; 
				4'b0001 : d <=  32'b00000000000000000000000000000110;
				4'b0010 : d <=  32'b00000000000000000000000000001100; 
				4'b0011 : d <=  32'b00000000000000000000000000000111; 
				4'b0100 : d <=  32'b00000000000000000000000000001111; 
				4'b0101 : d <=  32'b00000000000000000000000000100111; 
				4'b0110 : d <=  32'b00000000000000000000000001000111; 
				4'b0111 : d <=  32'b00000000000000000000000000101111;
				4'b1000 : d <=  32'b00000000000000000000000000100000;
				4'b1001 : d <=  32'b00000000000000000000000000100010;
				4'b1010 : d <=  32'b00000000000000000000000000100001;
				4'b1011 : d <=  32'b00000000000000000000000000100110;
				4'b1100 : d <=  32'b00000000000000000000000000111111;
				4'b1101 : d <=  32'b00000000000000000000000010001000;
				4'b1110 : d <=  32'b00000000000000000000000001100000;	
				4'b1111 : d <=  32'b00000000000000000000000001100001;	
							    
				default : d <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;	
			endcase//FIN case addr
			
			default : d <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
		endcase//FIN case en          
    end
endmodule
